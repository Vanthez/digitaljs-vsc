module a(
    input totally_identifiable_input, b,
    output c
);
and(c, totally_identifiable_input, b); 
endmodule
