module test(
    input a, b,
