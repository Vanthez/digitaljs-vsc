module test(
    input a, b,
    output c
);
and(c, a, b); 
endmodule
